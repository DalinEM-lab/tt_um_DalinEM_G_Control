VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_DalinEM_G_Control
  CLASS BLOCK ;
  FOREIGN tt_um_DalinEM_G_Control ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.000000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.000000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 259.387085 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 142.000 5.000 144.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 61.155 58.265 103.070 58.270 ;
        RECT 61.155 53.300 119.045 58.265 ;
        RECT 102.685 53.295 119.045 53.300 ;
      LAYER pwell ;
        RECT 64.495 47.590 131.675 47.605 ;
        RECT 61.305 44.025 131.675 47.590 ;
        RECT 61.305 44.010 64.585 44.025 ;
        RECT 67.690 42.025 106.115 44.025 ;
        RECT 118.810 35.025 125.285 44.025 ;
        RECT 61.065 16.125 122.175 31.455 ;
        RECT 126.060 16.110 133.990 41.930 ;
        RECT 134.415 16.105 136.425 26.925 ;
      LAYER li1 ;
        RECT 60.910 58.535 119.085 58.600 ;
        RECT 60.910 57.650 119.125 58.535 ;
        RECT 60.910 54.005 61.715 57.650 ;
        RECT 62.445 57.020 63.445 57.190 ;
        RECT 62.215 54.765 62.385 56.805 ;
        RECT 63.505 54.765 63.675 56.805 ;
        RECT 62.445 54.380 63.445 54.550 ;
        RECT 64.175 54.005 64.910 57.650 ;
        RECT 65.635 57.020 66.635 57.190 ;
        RECT 65.405 54.765 65.575 56.805 ;
        RECT 66.695 54.765 66.865 56.805 ;
        RECT 65.635 54.380 66.635 54.550 ;
        RECT 67.365 54.005 68.100 57.650 ;
        RECT 68.830 57.020 69.830 57.190 ;
        RECT 68.600 54.765 68.770 56.805 ;
        RECT 69.890 54.765 70.060 56.805 ;
        RECT 68.830 54.380 69.830 54.550 ;
        RECT 70.560 54.005 71.295 57.650 ;
        RECT 72.025 57.020 73.025 57.190 ;
        RECT 71.795 54.765 71.965 56.805 ;
        RECT 73.085 54.765 73.255 56.805 ;
        RECT 72.025 54.380 73.025 54.550 ;
        RECT 73.755 54.005 74.490 57.650 ;
        RECT 75.220 57.020 76.220 57.190 ;
        RECT 74.990 54.765 75.160 56.805 ;
        RECT 76.280 54.765 76.450 56.805 ;
        RECT 75.220 54.380 76.220 54.550 ;
        RECT 76.950 54.005 77.685 57.650 ;
        RECT 78.415 57.020 79.415 57.190 ;
        RECT 78.185 54.765 78.355 56.805 ;
        RECT 79.475 54.765 79.645 56.805 ;
        RECT 78.415 54.380 79.415 54.550 ;
        RECT 80.145 54.005 80.880 57.650 ;
        RECT 81.610 57.020 82.610 57.190 ;
        RECT 81.380 54.765 81.550 56.805 ;
        RECT 82.670 54.765 82.840 56.805 ;
        RECT 81.610 54.380 82.610 54.550 ;
        RECT 83.340 54.005 84.075 57.650 ;
        RECT 84.805 57.020 85.805 57.190 ;
        RECT 84.575 54.765 84.745 56.805 ;
        RECT 85.865 54.765 86.035 56.805 ;
        RECT 84.805 54.380 85.805 54.550 ;
        RECT 86.535 54.005 87.270 57.650 ;
        RECT 88.000 57.020 89.000 57.190 ;
        RECT 87.770 54.765 87.940 56.805 ;
        RECT 89.060 54.765 89.230 56.805 ;
        RECT 88.000 54.380 89.000 54.550 ;
        RECT 89.725 54.005 90.465 57.650 ;
        RECT 91.195 57.020 92.195 57.190 ;
        RECT 90.965 54.765 91.135 56.805 ;
        RECT 92.255 54.765 92.425 56.805 ;
        RECT 91.195 54.380 92.195 54.550 ;
        RECT 92.925 54.005 93.660 57.650 ;
        RECT 94.390 57.020 95.390 57.190 ;
        RECT 94.160 54.765 94.330 56.805 ;
        RECT 95.450 54.765 95.620 56.805 ;
        RECT 94.390 54.380 95.390 54.550 ;
        RECT 96.120 54.005 96.855 57.650 ;
        RECT 97.585 57.020 98.585 57.190 ;
        RECT 97.355 54.765 97.525 56.805 ;
        RECT 98.645 54.765 98.815 56.805 ;
        RECT 97.585 54.380 98.585 54.550 ;
        RECT 99.315 54.005 100.050 57.650 ;
        RECT 100.780 57.020 101.780 57.190 ;
        RECT 100.550 54.765 100.720 56.805 ;
        RECT 101.840 54.765 102.010 56.805 ;
        RECT 100.780 54.380 101.780 54.550 ;
        RECT 102.510 54.005 103.245 57.650 ;
        RECT 103.975 57.015 104.975 57.185 ;
        RECT 103.745 54.760 103.915 56.800 ;
        RECT 105.035 54.760 105.205 56.800 ;
        RECT 103.975 54.375 104.975 54.545 ;
        RECT 105.705 54.005 106.440 57.650 ;
        RECT 107.170 57.015 108.170 57.185 ;
        RECT 106.940 54.760 107.110 56.800 ;
        RECT 108.230 54.760 108.400 56.800 ;
        RECT 107.170 54.375 108.170 54.545 ;
        RECT 108.900 54.005 109.635 57.650 ;
        RECT 110.365 57.015 111.365 57.185 ;
        RECT 110.135 54.760 110.305 56.800 ;
        RECT 111.425 54.760 111.595 56.800 ;
        RECT 110.365 54.375 111.365 54.545 ;
        RECT 112.090 54.005 112.830 57.650 ;
        RECT 113.560 57.015 114.560 57.185 ;
        RECT 113.330 54.760 113.500 56.800 ;
        RECT 114.620 54.760 114.790 56.800 ;
        RECT 113.560 54.375 114.560 54.545 ;
        RECT 115.290 54.005 116.025 57.650 ;
        RECT 116.755 57.015 117.755 57.185 ;
        RECT 116.525 54.760 116.695 56.800 ;
        RECT 117.815 54.760 117.985 56.800 ;
        RECT 116.755 54.375 117.755 54.545 ;
        RECT 118.435 54.005 119.125 57.650 ;
        RECT 60.910 53.410 119.125 54.005 ;
        RECT 60.910 53.295 119.085 53.410 ;
        RECT 60.470 47.635 131.555 47.645 ;
        RECT 60.470 47.605 131.765 47.635 ;
        RECT 60.470 47.590 131.805 47.605 ;
        RECT 60.420 47.070 131.805 47.590 ;
        RECT 60.420 44.515 61.800 47.070 ;
        RECT 62.445 46.490 63.445 46.660 ;
        RECT 62.215 45.280 62.385 46.320 ;
        RECT 63.505 45.280 63.675 46.320 ;
        RECT 62.445 44.940 63.445 45.110 ;
        RECT 64.175 44.515 64.905 47.070 ;
        RECT 65.635 46.505 66.635 46.675 ;
        RECT 65.405 45.295 65.575 46.335 ;
        RECT 66.695 45.295 66.865 46.335 ;
        RECT 65.635 44.955 66.635 45.125 ;
        RECT 67.365 44.515 68.100 47.070 ;
        RECT 68.830 46.505 69.830 46.675 ;
        RECT 60.420 42.620 68.100 44.515 ;
        RECT 68.600 43.295 68.770 46.335 ;
        RECT 69.890 43.295 70.060 46.335 ;
        RECT 68.830 42.955 69.830 43.125 ;
        RECT 70.560 42.620 71.295 47.070 ;
        RECT 72.025 46.505 73.025 46.675 ;
        RECT 71.795 43.295 71.965 46.335 ;
        RECT 73.085 43.295 73.255 46.335 ;
        RECT 72.025 42.955 73.025 43.125 ;
        RECT 73.755 42.620 74.490 47.070 ;
        RECT 75.220 46.505 76.220 46.675 ;
        RECT 74.990 43.295 75.160 46.335 ;
        RECT 76.280 43.295 76.450 46.335 ;
        RECT 75.220 42.955 76.220 43.125 ;
        RECT 76.950 42.620 77.685 47.070 ;
        RECT 78.415 46.505 79.415 46.675 ;
        RECT 78.185 43.295 78.355 46.335 ;
        RECT 79.475 43.295 79.645 46.335 ;
        RECT 78.415 42.955 79.415 43.125 ;
        RECT 80.145 42.620 80.880 47.070 ;
        RECT 81.610 46.505 82.610 46.675 ;
        RECT 81.380 43.295 81.550 46.335 ;
        RECT 82.670 43.295 82.840 46.335 ;
        RECT 81.610 42.955 82.610 43.125 ;
        RECT 83.340 42.620 84.075 47.070 ;
        RECT 84.805 46.505 85.805 46.675 ;
        RECT 84.575 43.295 84.745 46.335 ;
        RECT 85.865 43.295 86.035 46.335 ;
        RECT 84.805 42.955 85.805 43.125 ;
        RECT 86.535 42.620 87.270 47.070 ;
        RECT 88.000 46.505 89.000 46.675 ;
        RECT 87.770 43.295 87.940 46.335 ;
        RECT 89.060 43.295 89.230 46.335 ;
        RECT 88.000 42.955 89.000 43.125 ;
        RECT 89.730 42.620 90.465 47.070 ;
        RECT 91.195 46.505 92.195 46.675 ;
        RECT 90.965 43.295 91.135 46.335 ;
        RECT 92.255 43.295 92.425 46.335 ;
        RECT 91.195 42.955 92.195 43.125 ;
        RECT 92.925 42.620 93.660 47.070 ;
        RECT 94.390 46.505 95.390 46.675 ;
        RECT 94.160 43.295 94.330 46.335 ;
        RECT 95.450 43.295 95.620 46.335 ;
        RECT 94.390 42.955 95.390 43.125 ;
        RECT 96.120 42.620 96.855 47.070 ;
        RECT 97.585 46.505 98.585 46.675 ;
        RECT 97.355 43.295 97.525 46.335 ;
        RECT 98.645 43.295 98.815 46.335 ;
        RECT 97.585 42.955 98.585 43.125 ;
        RECT 99.315 42.620 100.050 47.070 ;
        RECT 100.780 46.505 101.780 46.675 ;
        RECT 100.550 43.295 100.720 46.335 ;
        RECT 101.840 43.295 102.010 46.335 ;
        RECT 100.780 42.955 101.780 43.125 ;
        RECT 102.510 42.620 103.245 47.070 ;
        RECT 103.975 46.505 104.975 46.675 ;
        RECT 103.745 43.295 103.915 46.335 ;
        RECT 105.035 43.295 105.205 46.335 ;
        RECT 105.705 44.435 106.440 47.070 ;
        RECT 107.170 46.505 108.170 46.675 ;
        RECT 106.940 45.295 107.110 46.335 ;
        RECT 108.230 45.295 108.400 46.335 ;
        RECT 107.170 44.955 108.170 45.125 ;
        RECT 108.900 44.435 109.635 47.070 ;
        RECT 110.365 46.505 111.365 46.675 ;
        RECT 110.135 45.295 110.305 46.335 ;
        RECT 111.425 45.295 111.595 46.335 ;
        RECT 110.365 44.955 111.365 45.125 ;
        RECT 112.095 44.435 112.830 47.070 ;
        RECT 113.560 46.505 114.560 46.675 ;
        RECT 113.330 45.295 113.500 46.335 ;
        RECT 114.620 45.295 114.790 46.335 ;
        RECT 113.560 44.955 114.560 45.125 ;
        RECT 115.290 44.435 116.025 47.070 ;
        RECT 116.755 46.505 117.755 46.675 ;
        RECT 116.525 45.295 116.695 46.335 ;
        RECT 117.815 45.295 117.985 46.335 ;
        RECT 116.755 44.955 117.755 45.125 ;
        RECT 118.485 44.465 119.220 47.070 ;
        RECT 119.950 46.505 120.950 46.675 ;
        RECT 117.805 44.435 119.220 44.465 ;
        RECT 103.975 42.955 104.975 43.125 ;
        RECT 105.705 42.620 119.220 44.435 ;
        RECT 60.420 35.615 119.220 42.620 ;
        RECT 119.720 36.295 119.890 46.335 ;
        RECT 121.010 36.295 121.180 46.335 ;
        RECT 119.950 35.955 120.950 36.125 ;
        RECT 121.680 35.615 122.415 47.070 ;
        RECT 123.145 46.505 124.145 46.675 ;
        RECT 122.915 36.295 123.085 46.335 ;
        RECT 124.205 36.295 124.375 46.335 ;
        RECT 124.875 44.515 125.630 47.070 ;
        RECT 126.340 46.505 127.340 46.675 ;
        RECT 126.110 45.295 126.280 46.335 ;
        RECT 127.400 45.295 127.570 46.335 ;
        RECT 126.340 44.955 127.340 45.125 ;
        RECT 128.070 44.515 128.805 47.070 ;
        RECT 129.535 46.505 130.535 46.675 ;
        RECT 129.305 45.295 129.475 46.335 ;
        RECT 130.595 45.295 130.765 46.335 ;
        RECT 129.535 44.955 130.535 45.125 ;
        RECT 131.210 44.515 131.805 47.070 ;
        RECT 124.875 42.220 131.805 44.515 ;
        RECT 124.875 41.525 134.500 42.220 ;
        RECT 123.145 35.955 124.145 36.125 ;
        RECT 124.875 35.615 126.480 41.525 ;
        RECT 126.890 38.940 127.240 41.100 ;
        RECT 60.420 35.570 126.480 35.615 ;
        RECT 60.420 31.010 126.510 35.570 ;
        RECT 60.420 30.005 61.460 31.010 ;
        RECT 61.895 30.275 64.055 30.625 ;
        RECT 88.895 30.275 91.055 30.625 ;
        RECT 91.535 30.005 91.705 31.010 ;
        RECT 92.185 30.275 94.345 30.625 ;
        RECT 119.185 30.275 121.345 30.625 ;
        RECT 121.735 30.005 126.510 31.010 ;
        RECT 60.420 29.480 126.510 30.005 ;
        RECT 60.420 28.510 61.460 29.480 ;
        RECT 61.895 28.795 64.055 29.145 ;
        RECT 88.895 28.795 91.055 29.145 ;
        RECT 91.535 28.510 91.705 29.480 ;
        RECT 92.185 28.795 94.345 29.145 ;
        RECT 119.185 28.795 121.345 29.145 ;
        RECT 121.735 28.510 126.510 29.480 ;
        RECT 60.420 27.985 126.510 28.510 ;
        RECT 60.420 26.980 61.460 27.985 ;
        RECT 61.895 27.315 64.055 27.665 ;
        RECT 88.895 27.315 91.055 27.665 ;
        RECT 91.535 26.980 91.705 27.985 ;
        RECT 92.185 27.315 94.345 27.665 ;
        RECT 119.185 27.315 121.345 27.665 ;
        RECT 121.735 26.980 126.510 27.985 ;
        RECT 60.420 26.455 126.510 26.980 ;
        RECT 60.420 25.530 61.460 26.455 ;
        RECT 61.895 25.835 64.055 26.185 ;
        RECT 88.895 25.835 91.055 26.185 ;
        RECT 91.535 25.530 91.705 26.455 ;
        RECT 92.185 25.835 94.345 26.185 ;
        RECT 119.185 25.835 121.345 26.185 ;
        RECT 121.735 25.530 126.510 26.455 ;
        RECT 60.420 25.005 126.510 25.530 ;
        RECT 60.420 24.085 61.460 25.005 ;
        RECT 61.895 24.355 64.055 24.705 ;
        RECT 88.895 24.355 91.055 24.705 ;
        RECT 91.535 24.085 91.705 25.005 ;
        RECT 92.185 24.355 94.345 24.705 ;
        RECT 119.185 24.355 121.345 24.705 ;
        RECT 121.735 24.085 126.510 25.005 ;
        RECT 60.420 23.560 126.510 24.085 ;
        RECT 60.420 22.595 61.460 23.560 ;
        RECT 61.895 22.875 64.055 23.225 ;
        RECT 88.895 22.875 91.055 23.225 ;
        RECT 91.535 22.595 91.705 23.560 ;
        RECT 92.185 22.875 94.345 23.225 ;
        RECT 119.185 22.875 121.345 23.225 ;
        RECT 121.735 22.595 126.510 23.560 ;
        RECT 60.420 22.070 126.510 22.595 ;
        RECT 60.420 21.145 61.460 22.070 ;
        RECT 61.895 21.395 64.055 21.745 ;
        RECT 88.895 21.395 91.055 21.745 ;
        RECT 91.535 21.145 91.705 22.070 ;
        RECT 92.185 21.395 94.345 21.745 ;
        RECT 119.185 21.395 121.345 21.745 ;
        RECT 121.735 21.145 126.510 22.070 ;
        RECT 60.420 20.620 126.510 21.145 ;
        RECT 60.420 19.615 61.460 20.620 ;
        RECT 61.895 19.915 64.055 20.265 ;
        RECT 88.895 19.915 91.055 20.265 ;
        RECT 91.535 19.615 91.705 20.620 ;
        RECT 92.185 19.915 94.345 20.265 ;
        RECT 119.185 19.915 121.345 20.265 ;
        RECT 121.735 19.615 126.510 20.620 ;
        RECT 60.420 19.090 126.510 19.615 ;
        RECT 60.420 18.210 61.460 19.090 ;
        RECT 61.895 18.435 64.055 18.785 ;
        RECT 88.895 18.435 91.055 18.785 ;
        RECT 91.535 18.210 91.705 19.090 ;
        RECT 92.185 18.435 94.345 18.785 ;
        RECT 119.185 18.435 121.345 18.785 ;
        RECT 121.735 18.210 126.510 19.090 ;
        RECT 60.420 17.685 126.510 18.210 ;
        RECT 60.420 16.610 61.460 17.685 ;
        RECT 61.895 16.955 64.055 17.305 ;
        RECT 88.895 16.955 91.055 17.305 ;
        RECT 91.535 16.610 91.705 17.685 ;
        RECT 92.185 16.955 94.345 17.305 ;
        RECT 119.185 16.955 121.345 17.305 ;
        RECT 121.735 16.610 126.510 17.685 ;
        RECT 126.890 16.940 127.240 19.100 ;
        RECT 60.400 16.545 126.510 16.610 ;
        RECT 127.595 16.545 128.090 41.525 ;
        RECT 128.370 38.940 128.720 41.100 ;
        RECT 128.370 16.940 128.720 19.100 ;
        RECT 129.045 16.545 129.540 41.525 ;
        RECT 129.850 38.940 130.200 41.100 ;
        RECT 129.850 16.940 130.200 19.100 ;
        RECT 130.540 16.545 131.035 41.525 ;
        RECT 131.330 38.940 131.680 41.100 ;
        RECT 131.330 16.940 131.680 19.100 ;
        RECT 132.030 16.545 132.525 41.525 ;
        RECT 132.810 38.940 133.160 41.100 ;
        RECT 133.570 27.025 134.450 41.525 ;
        RECT 137.590 27.185 137.850 28.680 ;
        RECT 133.570 26.425 136.790 27.025 ;
        RECT 137.225 26.900 138.225 27.185 ;
        RECT 132.810 16.940 133.160 19.100 ;
        RECT 133.570 16.545 134.780 26.425 ;
        RECT 135.245 23.935 135.595 26.095 ;
        RECT 135.245 16.935 135.595 19.095 ;
        RECT 60.400 16.490 134.780 16.545 ;
        RECT 136.060 16.495 136.740 26.425 ;
        RECT 137.225 16.615 138.225 16.900 ;
        RECT 135.930 16.490 136.760 16.495 ;
        RECT 60.400 15.665 136.760 16.490 ;
        RECT 137.580 15.720 137.990 16.615 ;
        RECT 125.730 15.615 136.760 15.665 ;
      LAYER met1 ;
        RECT 60.930 58.500 61.610 58.540 ;
        RECT 118.475 58.535 119.155 58.595 ;
        RECT 118.455 58.500 119.175 58.535 ;
        RECT 60.930 58.480 119.175 58.500 ;
        RECT 60.910 57.725 119.175 58.480 ;
        RECT 60.910 53.950 61.630 57.725 ;
        RECT 62.465 56.990 63.425 57.220 ;
        RECT 62.185 56.725 62.415 56.785 ;
        RECT 62.120 56.325 62.480 56.725 ;
        RECT 62.185 54.785 62.415 56.325 ;
        RECT 63.475 55.245 63.705 56.785 ;
        RECT 63.410 54.845 63.770 55.245 ;
        RECT 63.475 54.785 63.705 54.845 ;
        RECT 62.475 54.580 62.975 54.595 ;
        RECT 62.465 54.350 63.425 54.580 ;
        RECT 62.475 54.335 62.975 54.350 ;
        RECT 64.215 53.950 64.860 57.725 ;
        RECT 65.655 56.990 66.615 57.220 ;
        RECT 65.375 56.725 65.605 56.785 ;
        RECT 65.310 56.325 65.670 56.725 ;
        RECT 65.375 54.785 65.605 56.325 ;
        RECT 66.665 55.245 66.895 56.785 ;
        RECT 66.600 54.845 66.960 55.245 ;
        RECT 66.665 54.785 66.895 54.845 ;
        RECT 65.665 54.580 66.165 54.595 ;
        RECT 65.655 54.350 66.615 54.580 ;
        RECT 65.665 54.335 66.165 54.350 ;
        RECT 67.425 53.950 68.070 57.725 ;
        RECT 68.850 56.990 69.810 57.220 ;
        RECT 68.570 55.245 68.800 56.785 ;
        RECT 69.860 56.725 70.090 56.785 ;
        RECT 69.795 56.325 70.155 56.725 ;
        RECT 68.505 54.845 68.865 55.245 ;
        RECT 68.570 54.785 68.800 54.845 ;
        RECT 69.860 54.785 70.090 56.325 ;
        RECT 69.300 54.580 69.800 54.590 ;
        RECT 68.850 54.350 69.810 54.580 ;
        RECT 69.300 54.330 69.800 54.350 ;
        RECT 70.635 53.950 71.280 57.725 ;
        RECT 72.045 56.990 73.005 57.220 ;
        RECT 71.765 55.245 71.995 56.785 ;
        RECT 73.055 56.725 73.285 56.785 ;
        RECT 72.990 56.325 73.350 56.725 ;
        RECT 71.700 54.845 72.060 55.245 ;
        RECT 71.765 54.785 71.995 54.845 ;
        RECT 73.055 54.785 73.285 56.325 ;
        RECT 72.495 54.580 72.995 54.595 ;
        RECT 72.045 54.350 73.005 54.580 ;
        RECT 72.495 54.335 72.995 54.350 ;
        RECT 73.795 53.950 74.440 57.725 ;
        RECT 75.240 56.990 76.200 57.220 ;
        RECT 74.960 55.245 75.190 56.785 ;
        RECT 76.250 56.725 76.480 56.785 ;
        RECT 76.185 56.325 76.545 56.725 ;
        RECT 74.895 54.845 75.255 55.245 ;
        RECT 74.960 54.785 75.190 54.845 ;
        RECT 76.250 54.785 76.480 56.325 ;
        RECT 75.690 54.580 76.190 54.595 ;
        RECT 75.240 54.350 76.200 54.580 ;
        RECT 75.690 54.335 76.190 54.350 ;
        RECT 77.000 53.950 77.645 57.725 ;
        RECT 78.435 56.990 79.395 57.220 ;
        RECT 78.155 55.245 78.385 56.785 ;
        RECT 79.445 56.725 79.675 56.785 ;
        RECT 79.380 56.325 79.740 56.725 ;
        RECT 78.090 54.845 78.450 55.245 ;
        RECT 78.155 54.785 78.385 54.845 ;
        RECT 79.445 54.785 79.675 56.325 ;
        RECT 78.885 54.580 79.385 54.595 ;
        RECT 78.435 54.350 79.395 54.580 ;
        RECT 78.885 54.335 79.385 54.350 ;
        RECT 80.205 53.950 80.850 57.725 ;
        RECT 81.630 56.990 82.590 57.220 ;
        RECT 81.350 55.245 81.580 56.785 ;
        RECT 82.640 56.725 82.870 56.785 ;
        RECT 82.575 56.325 82.935 56.725 ;
        RECT 81.285 54.845 81.645 55.245 ;
        RECT 81.350 54.785 81.580 54.845 ;
        RECT 82.640 54.785 82.870 56.325 ;
        RECT 82.080 54.580 82.580 54.595 ;
        RECT 81.630 54.350 82.590 54.580 ;
        RECT 82.080 54.335 82.580 54.350 ;
        RECT 83.430 53.950 84.075 57.725 ;
        RECT 84.825 56.990 85.785 57.220 ;
        RECT 84.545 55.245 84.775 56.785 ;
        RECT 85.835 56.725 86.065 56.785 ;
        RECT 85.770 56.325 86.130 56.725 ;
        RECT 84.480 54.845 84.840 55.245 ;
        RECT 84.545 54.785 84.775 54.845 ;
        RECT 85.835 54.785 86.065 56.325 ;
        RECT 85.275 54.580 85.775 54.595 ;
        RECT 84.825 54.350 85.785 54.580 ;
        RECT 85.275 54.335 85.775 54.350 ;
        RECT 85.320 53.950 85.905 53.955 ;
        RECT 86.545 53.950 87.190 57.725 ;
        RECT 88.020 56.990 88.980 57.220 ;
        RECT 87.740 55.245 87.970 56.785 ;
        RECT 89.030 56.725 89.260 56.785 ;
        RECT 88.965 56.325 89.325 56.725 ;
        RECT 87.675 54.845 88.035 55.245 ;
        RECT 87.740 54.785 87.970 54.845 ;
        RECT 89.030 54.785 89.260 56.325 ;
        RECT 88.470 54.580 88.970 54.595 ;
        RECT 88.020 54.350 88.980 54.580 ;
        RECT 88.470 54.335 88.970 54.350 ;
        RECT 89.795 53.950 90.440 57.725 ;
        RECT 91.215 56.990 92.175 57.220 ;
        RECT 90.935 55.245 91.165 56.785 ;
        RECT 92.225 56.725 92.455 56.785 ;
        RECT 92.160 56.325 92.520 56.725 ;
        RECT 90.870 54.845 91.230 55.245 ;
        RECT 90.935 54.785 91.165 54.845 ;
        RECT 92.225 54.785 92.455 56.325 ;
        RECT 91.665 54.580 92.165 54.595 ;
        RECT 91.215 54.350 92.175 54.580 ;
        RECT 91.665 54.335 92.165 54.350 ;
        RECT 92.975 53.950 93.620 57.725 ;
        RECT 94.410 56.990 95.370 57.220 ;
        RECT 94.130 55.245 94.360 56.785 ;
        RECT 95.420 56.725 95.650 56.785 ;
        RECT 95.355 56.325 95.715 56.725 ;
        RECT 94.065 54.845 94.425 55.245 ;
        RECT 94.130 54.785 94.360 54.845 ;
        RECT 95.420 54.785 95.650 56.325 ;
        RECT 94.860 54.580 95.360 54.595 ;
        RECT 94.410 54.350 95.370 54.580 ;
        RECT 94.860 54.335 95.360 54.350 ;
        RECT 96.180 53.950 96.825 57.725 ;
        RECT 97.605 56.990 98.565 57.220 ;
        RECT 97.325 55.245 97.555 56.785 ;
        RECT 98.615 56.725 98.845 56.785 ;
        RECT 98.550 56.325 98.910 56.725 ;
        RECT 97.260 54.845 97.620 55.245 ;
        RECT 97.325 54.785 97.555 54.845 ;
        RECT 98.615 54.785 98.845 56.325 ;
        RECT 98.055 54.580 98.555 54.595 ;
        RECT 97.605 54.350 98.565 54.580 ;
        RECT 98.055 54.335 98.555 54.350 ;
        RECT 99.340 53.950 99.985 57.725 ;
        RECT 100.800 56.990 101.760 57.220 ;
        RECT 100.520 55.245 100.750 56.785 ;
        RECT 101.810 56.725 102.040 56.785 ;
        RECT 101.745 56.325 102.105 56.725 ;
        RECT 100.455 54.845 100.815 55.245 ;
        RECT 100.520 54.785 100.750 54.845 ;
        RECT 101.810 54.785 102.040 56.325 ;
        RECT 101.250 54.580 101.750 54.595 ;
        RECT 100.800 54.350 101.760 54.580 ;
        RECT 101.250 54.335 101.750 54.350 ;
        RECT 102.565 53.950 103.210 57.725 ;
        RECT 103.995 56.985 104.955 57.215 ;
        RECT 103.715 55.240 103.945 56.780 ;
        RECT 105.005 56.720 105.235 56.780 ;
        RECT 104.940 56.320 105.300 56.720 ;
        RECT 103.650 54.840 104.010 55.240 ;
        RECT 103.715 54.780 103.945 54.840 ;
        RECT 105.005 54.780 105.235 56.320 ;
        RECT 104.445 54.575 104.945 54.590 ;
        RECT 103.995 54.345 104.955 54.575 ;
        RECT 104.445 54.330 104.945 54.345 ;
        RECT 105.750 53.950 106.395 57.725 ;
        RECT 107.190 56.985 108.150 57.215 ;
        RECT 106.910 56.720 107.140 56.780 ;
        RECT 106.845 56.320 107.205 56.720 ;
        RECT 106.910 54.780 107.140 56.320 ;
        RECT 108.200 55.240 108.430 56.780 ;
        RECT 108.135 54.840 108.495 55.240 ;
        RECT 108.200 54.780 108.430 54.840 ;
        RECT 107.200 54.575 107.700 54.590 ;
        RECT 107.190 54.345 108.150 54.575 ;
        RECT 107.200 54.330 107.700 54.345 ;
        RECT 108.975 53.950 109.620 57.725 ;
        RECT 110.385 56.985 111.345 57.215 ;
        RECT 110.105 56.720 110.335 56.780 ;
        RECT 110.040 56.320 110.400 56.720 ;
        RECT 110.105 54.780 110.335 56.320 ;
        RECT 111.395 55.240 111.625 56.780 ;
        RECT 111.330 54.840 111.690 55.240 ;
        RECT 111.395 54.780 111.625 54.840 ;
        RECT 110.395 54.575 110.895 54.590 ;
        RECT 110.385 54.345 111.345 54.575 ;
        RECT 110.395 54.330 110.895 54.345 ;
        RECT 112.180 53.950 112.825 57.725 ;
        RECT 113.580 56.985 114.540 57.215 ;
        RECT 113.300 56.720 113.530 56.780 ;
        RECT 113.235 56.320 113.595 56.720 ;
        RECT 113.300 54.780 113.530 56.320 ;
        RECT 114.590 55.240 114.820 56.780 ;
        RECT 114.525 54.840 114.885 55.240 ;
        RECT 114.590 54.780 114.820 54.840 ;
        RECT 113.590 54.575 114.090 54.590 ;
        RECT 113.580 54.345 114.540 54.575 ;
        RECT 113.590 54.330 114.090 54.345 ;
        RECT 115.360 53.950 116.005 57.725 ;
        RECT 116.775 56.985 117.735 57.215 ;
        RECT 116.495 56.720 116.725 56.780 ;
        RECT 116.430 56.320 116.790 56.720 ;
        RECT 116.495 54.780 116.725 56.320 ;
        RECT 117.785 55.240 118.015 56.780 ;
        RECT 117.720 54.840 118.080 55.240 ;
        RECT 117.785 54.780 118.015 54.840 ;
        RECT 116.785 54.575 117.285 54.590 ;
        RECT 116.775 54.345 117.735 54.575 ;
        RECT 116.785 54.330 117.285 54.345 ;
        RECT 118.455 53.950 119.175 57.725 ;
        RECT 60.910 53.410 119.175 53.950 ;
        RECT 60.910 53.355 119.155 53.410 ;
        RECT 60.930 53.350 119.155 53.355 ;
        RECT 60.930 53.300 119.030 53.350 ;
        RECT 60.930 53.295 61.610 53.300 ;
        RECT 56.990 49.325 60.035 49.540 ;
        RECT 56.990 49.025 66.055 49.325 ;
        RECT 56.990 48.640 60.035 49.025 ;
        RECT 56.990 39.105 57.890 48.640 ;
        RECT 131.180 47.620 131.835 47.665 ;
        RECT 60.360 47.375 131.835 47.620 ;
        RECT 60.370 47.110 131.835 47.375 ;
        RECT 60.370 44.545 61.310 47.110 ;
        RECT 65.665 46.705 66.165 46.720 ;
        RECT 69.300 46.705 69.800 46.720 ;
        RECT 72.495 46.705 72.995 46.720 ;
        RECT 75.690 46.705 76.190 46.720 ;
        RECT 78.885 46.705 79.385 46.720 ;
        RECT 82.080 46.705 82.580 46.720 ;
        RECT 85.275 46.705 85.775 46.720 ;
        RECT 88.470 46.705 88.970 46.720 ;
        RECT 91.665 46.705 92.165 46.720 ;
        RECT 94.860 46.705 95.360 46.720 ;
        RECT 98.055 46.705 98.555 46.720 ;
        RECT 101.250 46.705 101.750 46.720 ;
        RECT 104.445 46.705 104.945 46.720 ;
        RECT 107.200 46.705 107.700 46.720 ;
        RECT 110.395 46.705 110.895 46.720 ;
        RECT 113.590 46.705 114.090 46.720 ;
        RECT 116.785 46.705 117.285 46.720 ;
        RECT 119.980 46.705 120.480 46.720 ;
        RECT 62.475 46.690 62.975 46.705 ;
        RECT 62.465 46.460 63.425 46.690 ;
        RECT 65.655 46.475 66.615 46.705 ;
        RECT 68.850 46.475 69.810 46.705 ;
        RECT 72.045 46.475 73.005 46.705 ;
        RECT 75.240 46.475 76.200 46.705 ;
        RECT 78.435 46.475 79.395 46.705 ;
        RECT 81.630 46.475 82.590 46.705 ;
        RECT 84.825 46.475 85.785 46.705 ;
        RECT 88.020 46.475 88.980 46.705 ;
        RECT 91.215 46.475 92.175 46.705 ;
        RECT 94.410 46.475 95.370 46.705 ;
        RECT 97.605 46.475 98.565 46.705 ;
        RECT 100.800 46.475 101.760 46.705 ;
        RECT 103.995 46.475 104.955 46.705 ;
        RECT 107.190 46.475 108.150 46.705 ;
        RECT 110.385 46.475 111.345 46.705 ;
        RECT 113.580 46.475 114.540 46.705 ;
        RECT 116.775 46.475 117.735 46.705 ;
        RECT 119.970 46.475 120.930 46.705 ;
        RECT 65.665 46.460 66.165 46.475 ;
        RECT 69.300 46.460 69.800 46.475 ;
        RECT 72.495 46.460 72.995 46.475 ;
        RECT 75.690 46.460 76.190 46.475 ;
        RECT 78.885 46.460 79.385 46.475 ;
        RECT 82.080 46.460 82.580 46.475 ;
        RECT 85.275 46.460 85.775 46.475 ;
        RECT 88.470 46.460 88.970 46.475 ;
        RECT 91.665 46.460 92.165 46.475 ;
        RECT 94.860 46.460 95.360 46.475 ;
        RECT 98.055 46.460 98.555 46.475 ;
        RECT 101.250 46.460 101.750 46.475 ;
        RECT 104.445 46.460 104.945 46.475 ;
        RECT 107.200 46.460 107.700 46.475 ;
        RECT 110.395 46.460 110.895 46.475 ;
        RECT 113.590 46.460 114.090 46.475 ;
        RECT 116.785 46.460 117.285 46.475 ;
        RECT 119.980 46.460 120.480 46.475 ;
        RECT 62.475 46.445 62.975 46.460 ;
        RECT 62.185 45.760 62.415 46.300 ;
        RECT 63.475 46.240 63.705 46.300 ;
        RECT 63.410 45.840 63.770 46.240 ;
        RECT 62.120 45.360 62.480 45.760 ;
        RECT 62.185 45.300 62.415 45.360 ;
        RECT 63.475 45.300 63.705 45.840 ;
        RECT 65.375 45.775 65.605 46.315 ;
        RECT 66.665 46.255 66.895 46.315 ;
        RECT 68.570 46.255 68.800 46.315 ;
        RECT 66.600 45.855 66.960 46.255 ;
        RECT 68.505 45.855 68.865 46.255 ;
        RECT 65.310 45.375 65.670 45.775 ;
        RECT 65.375 45.315 65.605 45.375 ;
        RECT 66.665 45.315 66.895 45.855 ;
        RECT 62.465 44.910 63.425 45.140 ;
        RECT 65.655 44.925 66.615 45.155 ;
        RECT 60.370 44.460 68.085 44.545 ;
        RECT 60.370 43.320 68.100 44.460 ;
        RECT 60.390 43.290 68.100 43.320 ;
        RECT 68.570 43.315 68.800 45.855 ;
        RECT 69.860 43.775 70.090 46.315 ;
        RECT 71.765 43.775 71.995 46.315 ;
        RECT 73.055 43.775 73.285 46.315 ;
        RECT 74.960 43.775 75.190 46.315 ;
        RECT 76.250 43.775 76.480 46.315 ;
        RECT 78.155 46.255 78.385 46.315 ;
        RECT 78.090 45.855 78.450 46.255 ;
        RECT 69.795 43.375 70.155 43.775 ;
        RECT 71.700 43.375 72.060 43.775 ;
        RECT 72.990 43.375 73.350 43.775 ;
        RECT 74.895 43.375 75.255 43.775 ;
        RECT 76.185 43.375 76.545 43.775 ;
        RECT 69.860 43.315 70.090 43.375 ;
        RECT 71.765 43.315 71.995 43.375 ;
        RECT 73.055 43.315 73.285 43.375 ;
        RECT 74.960 43.315 75.190 43.375 ;
        RECT 76.250 43.315 76.480 43.375 ;
        RECT 78.155 43.315 78.385 45.855 ;
        RECT 79.445 43.775 79.675 46.315 ;
        RECT 81.350 43.775 81.580 46.315 ;
        RECT 82.640 43.775 82.870 46.315 ;
        RECT 84.545 43.775 84.775 46.315 ;
        RECT 85.835 43.775 86.065 46.315 ;
        RECT 87.740 46.255 87.970 46.315 ;
        RECT 87.675 45.855 88.035 46.255 ;
        RECT 79.380 43.375 79.740 43.775 ;
        RECT 81.285 43.375 81.645 43.775 ;
        RECT 82.575 43.375 82.935 43.775 ;
        RECT 84.480 43.375 84.840 43.775 ;
        RECT 85.770 43.375 86.130 43.775 ;
        RECT 79.445 43.315 79.675 43.375 ;
        RECT 81.350 43.315 81.580 43.375 ;
        RECT 82.640 43.315 82.870 43.375 ;
        RECT 84.545 43.315 84.775 43.375 ;
        RECT 85.835 43.315 86.065 43.375 ;
        RECT 87.740 43.315 87.970 45.855 ;
        RECT 89.030 43.775 89.260 46.315 ;
        RECT 90.935 43.775 91.165 46.315 ;
        RECT 92.225 43.775 92.455 46.315 ;
        RECT 94.130 43.775 94.360 46.315 ;
        RECT 95.420 43.775 95.650 46.315 ;
        RECT 97.325 46.255 97.555 46.315 ;
        RECT 97.260 45.855 97.620 46.255 ;
        RECT 88.965 43.375 89.325 43.775 ;
        RECT 90.870 43.375 91.230 43.775 ;
        RECT 92.160 43.375 92.520 43.775 ;
        RECT 94.065 43.375 94.425 43.775 ;
        RECT 95.355 43.375 95.715 43.775 ;
        RECT 89.030 43.315 89.260 43.375 ;
        RECT 90.935 43.315 91.165 43.375 ;
        RECT 92.225 43.315 92.455 43.375 ;
        RECT 94.130 43.315 94.360 43.375 ;
        RECT 95.420 43.315 95.650 43.375 ;
        RECT 97.325 43.315 97.555 45.855 ;
        RECT 98.615 43.775 98.845 46.315 ;
        RECT 100.520 43.775 100.750 46.315 ;
        RECT 101.810 43.775 102.040 46.315 ;
        RECT 103.715 43.775 103.945 46.315 ;
        RECT 105.005 43.775 105.235 46.315 ;
        RECT 106.910 45.775 107.140 46.315 ;
        RECT 108.200 46.255 108.430 46.315 ;
        RECT 108.135 45.855 108.495 46.255 ;
        RECT 106.845 45.375 107.205 45.775 ;
        RECT 106.910 45.315 107.140 45.375 ;
        RECT 108.200 45.315 108.430 45.855 ;
        RECT 110.105 45.775 110.335 46.315 ;
        RECT 111.395 46.255 111.625 46.315 ;
        RECT 111.330 45.855 111.690 46.255 ;
        RECT 110.040 45.375 110.400 45.775 ;
        RECT 110.105 45.315 110.335 45.375 ;
        RECT 111.395 45.315 111.625 45.855 ;
        RECT 113.300 45.775 113.530 46.315 ;
        RECT 114.590 46.255 114.820 46.315 ;
        RECT 114.525 45.855 114.885 46.255 ;
        RECT 113.235 45.375 113.595 45.775 ;
        RECT 113.300 45.315 113.530 45.375 ;
        RECT 114.590 45.315 114.820 45.855 ;
        RECT 116.495 45.775 116.725 46.315 ;
        RECT 117.785 46.255 118.015 46.315 ;
        RECT 117.720 45.855 118.080 46.255 ;
        RECT 116.430 45.375 116.790 45.775 ;
        RECT 116.495 45.315 116.725 45.375 ;
        RECT 117.785 45.315 118.015 45.855 ;
        RECT 107.190 44.925 108.150 45.155 ;
        RECT 110.385 44.925 111.345 45.155 ;
        RECT 113.580 44.925 114.540 45.155 ;
        RECT 116.775 44.925 117.735 45.155 ;
        RECT 105.815 44.470 107.120 44.475 ;
        RECT 117.775 44.470 119.230 44.525 ;
        RECT 105.815 44.425 119.250 44.470 ;
        RECT 98.550 43.375 98.910 43.775 ;
        RECT 100.455 43.375 100.815 43.775 ;
        RECT 101.745 43.375 102.105 43.775 ;
        RECT 103.650 43.375 104.010 43.775 ;
        RECT 104.940 43.375 105.300 43.775 ;
        RECT 98.615 43.315 98.845 43.375 ;
        RECT 100.520 43.315 100.750 43.375 ;
        RECT 101.810 43.315 102.040 43.375 ;
        RECT 103.715 43.315 103.945 43.375 ;
        RECT 105.005 43.315 105.235 43.375 ;
        RECT 56.960 38.205 57.920 39.105 ;
        RECT 60.390 31.935 61.285 43.290 ;
        RECT 66.715 42.650 68.100 43.290 ;
        RECT 105.700 43.290 119.250 44.425 ;
        RECT 68.850 42.925 69.810 43.155 ;
        RECT 72.045 42.925 73.005 43.155 ;
        RECT 75.240 42.925 76.200 43.155 ;
        RECT 78.435 42.925 79.395 43.155 ;
        RECT 81.630 42.925 82.590 43.155 ;
        RECT 84.825 42.925 85.785 43.155 ;
        RECT 88.020 42.925 88.980 43.155 ;
        RECT 91.215 42.925 92.175 43.155 ;
        RECT 94.410 42.925 95.370 43.155 ;
        RECT 97.605 42.925 98.565 43.155 ;
        RECT 100.800 42.925 101.760 43.155 ;
        RECT 103.995 42.925 104.955 43.155 ;
        RECT 105.700 42.650 107.120 43.290 ;
        RECT 66.715 41.645 107.120 42.650 ;
        RECT 66.715 41.600 68.100 41.645 ;
        RECT 105.815 41.565 107.120 41.645 ;
        RECT 117.775 35.625 119.250 43.290 ;
        RECT 119.690 41.375 119.920 46.315 ;
        RECT 120.980 41.375 121.210 46.315 ;
        RECT 119.625 36.375 119.985 41.375 ;
        RECT 120.915 36.375 121.275 41.375 ;
        RECT 119.690 36.315 119.920 36.375 ;
        RECT 120.980 36.315 121.210 36.375 ;
        RECT 119.970 35.925 120.930 36.155 ;
        RECT 121.760 35.625 122.275 47.110 ;
        RECT 123.175 46.705 123.675 46.720 ;
        RECT 123.165 46.475 124.125 46.705 ;
        RECT 123.175 46.460 123.675 46.475 ;
        RECT 122.885 41.375 123.115 46.315 ;
        RECT 124.175 41.375 124.405 46.315 ;
        RECT 124.850 44.545 125.660 47.110 ;
        RECT 126.370 46.705 126.870 46.720 ;
        RECT 126.360 46.475 127.320 46.705 ;
        RECT 126.370 46.460 126.870 46.475 ;
        RECT 126.080 45.875 126.310 46.315 ;
        RECT 127.370 45.875 127.600 46.315 ;
        RECT 126.015 45.375 126.375 45.875 ;
        RECT 127.305 45.375 127.665 45.875 ;
        RECT 126.080 45.315 126.310 45.375 ;
        RECT 127.370 45.315 127.600 45.375 ;
        RECT 126.360 44.925 127.320 45.155 ;
        RECT 128.105 44.545 128.785 47.110 ;
        RECT 129.565 46.705 130.065 46.720 ;
        RECT 129.555 46.475 130.515 46.705 ;
        RECT 129.565 46.460 130.065 46.475 ;
        RECT 129.275 45.875 129.505 46.315 ;
        RECT 130.565 45.875 130.795 46.315 ;
        RECT 129.210 45.375 129.570 45.875 ;
        RECT 130.500 45.375 130.860 45.875 ;
        RECT 129.275 45.315 129.505 45.375 ;
        RECT 130.565 45.315 130.795 45.375 ;
        RECT 129.555 44.925 130.515 45.155 ;
        RECT 131.180 44.545 131.835 47.110 ;
        RECT 124.850 42.250 131.865 44.545 ;
        RECT 124.850 41.495 134.560 42.250 ;
        RECT 122.820 36.375 123.180 41.375 ;
        RECT 124.110 36.375 124.470 41.375 ;
        RECT 122.885 36.315 123.115 36.375 ;
        RECT 124.175 36.315 124.405 36.375 ;
        RECT 123.165 35.925 124.125 36.155 ;
        RECT 124.850 35.625 126.510 41.495 ;
        RECT 126.940 41.010 127.190 41.070 ;
        RECT 126.885 40.010 127.245 41.010 ;
        RECT 126.940 38.965 127.190 40.010 ;
        RECT 117.775 34.520 126.535 35.625 ;
        RECT 117.775 32.015 126.485 34.520 ;
        RECT 117.775 31.935 126.505 32.015 ;
        RECT 60.390 30.980 126.505 31.935 ;
        RECT 60.390 29.955 61.285 30.980 ;
        RECT 61.935 30.575 63.035 30.580 ;
        RECT 89.915 30.575 91.015 30.580 ;
        RECT 92.225 30.575 93.325 30.580 ;
        RECT 120.205 30.575 121.305 30.580 ;
        RECT 61.925 30.325 64.030 30.575 ;
        RECT 88.920 30.325 91.025 30.575 ;
        RECT 92.215 30.325 94.320 30.575 ;
        RECT 119.210 30.325 121.315 30.575 ;
        RECT 61.935 30.320 63.035 30.325 ;
        RECT 89.915 30.320 91.015 30.325 ;
        RECT 92.225 30.320 93.325 30.325 ;
        RECT 120.205 30.320 121.305 30.325 ;
        RECT 121.760 29.955 126.505 30.980 ;
        RECT 60.390 29.565 126.505 29.955 ;
        RECT 60.390 28.465 61.285 29.565 ;
        RECT 61.935 29.095 63.035 29.100 ;
        RECT 89.915 29.095 91.015 29.100 ;
        RECT 92.225 29.095 93.325 29.100 ;
        RECT 120.205 29.095 121.305 29.100 ;
        RECT 61.925 28.845 64.030 29.095 ;
        RECT 88.920 28.845 91.025 29.095 ;
        RECT 92.215 28.845 94.320 29.095 ;
        RECT 119.210 28.845 121.315 29.095 ;
        RECT 61.935 28.840 63.035 28.845 ;
        RECT 89.915 28.840 91.015 28.845 ;
        RECT 92.225 28.840 93.325 28.845 ;
        RECT 120.205 28.840 121.305 28.845 ;
        RECT 121.760 28.465 126.505 29.565 ;
        RECT 60.390 28.075 126.505 28.465 ;
        RECT 60.390 26.890 61.285 28.075 ;
        RECT 61.935 27.615 63.035 27.620 ;
        RECT 89.915 27.615 91.015 27.620 ;
        RECT 92.225 27.615 93.325 27.620 ;
        RECT 120.205 27.615 121.305 27.620 ;
        RECT 61.925 27.365 64.030 27.615 ;
        RECT 88.920 27.365 91.025 27.615 ;
        RECT 92.215 27.365 94.320 27.615 ;
        RECT 119.210 27.365 121.315 27.615 ;
        RECT 61.935 27.360 63.035 27.365 ;
        RECT 89.915 27.360 91.015 27.365 ;
        RECT 92.225 27.360 93.325 27.365 ;
        RECT 120.205 27.360 121.305 27.365 ;
        RECT 121.760 26.890 126.505 28.075 ;
        RECT 60.390 26.500 126.505 26.890 ;
        RECT 60.390 25.440 61.285 26.500 ;
        RECT 61.935 26.135 63.035 26.140 ;
        RECT 89.915 26.135 91.015 26.140 ;
        RECT 92.225 26.135 93.325 26.140 ;
        RECT 120.205 26.135 121.305 26.140 ;
        RECT 61.925 25.885 64.030 26.135 ;
        RECT 88.920 25.885 91.025 26.135 ;
        RECT 92.215 25.885 94.320 26.135 ;
        RECT 119.210 25.885 121.315 26.135 ;
        RECT 61.935 25.880 63.035 25.885 ;
        RECT 89.915 25.880 91.015 25.885 ;
        RECT 92.225 25.880 93.325 25.885 ;
        RECT 120.205 25.880 121.305 25.885 ;
        RECT 121.760 25.440 126.505 26.500 ;
        RECT 60.390 25.050 126.505 25.440 ;
        RECT 60.390 23.990 61.285 25.050 ;
        RECT 61.935 24.655 63.035 24.660 ;
        RECT 89.915 24.655 91.015 24.660 ;
        RECT 92.225 24.655 93.325 24.660 ;
        RECT 120.205 24.655 121.305 24.660 ;
        RECT 61.925 24.405 64.030 24.655 ;
        RECT 88.920 24.405 91.025 24.655 ;
        RECT 92.215 24.405 94.320 24.655 ;
        RECT 119.210 24.405 121.315 24.655 ;
        RECT 61.935 24.400 63.035 24.405 ;
        RECT 89.915 24.400 91.015 24.405 ;
        RECT 92.225 24.400 93.325 24.405 ;
        RECT 120.205 24.400 121.305 24.405 ;
        RECT 121.760 23.990 126.505 25.050 ;
        RECT 60.390 23.600 126.505 23.990 ;
        RECT 60.390 22.545 61.285 23.600 ;
        RECT 61.935 23.175 63.035 23.180 ;
        RECT 89.915 23.175 91.015 23.180 ;
        RECT 92.225 23.175 93.325 23.180 ;
        RECT 120.205 23.175 121.305 23.180 ;
        RECT 61.925 22.925 64.030 23.175 ;
        RECT 88.920 22.925 91.025 23.175 ;
        RECT 92.215 22.925 94.320 23.175 ;
        RECT 119.210 22.925 121.315 23.175 ;
        RECT 61.935 22.920 63.035 22.925 ;
        RECT 89.915 22.920 91.015 22.925 ;
        RECT 92.225 22.920 93.325 22.925 ;
        RECT 120.205 22.920 121.305 22.925 ;
        RECT 121.760 22.545 126.505 23.600 ;
        RECT 60.390 22.155 126.505 22.545 ;
        RECT 60.390 21.050 61.285 22.155 ;
        RECT 61.935 21.695 63.035 21.700 ;
        RECT 89.915 21.695 91.015 21.700 ;
        RECT 92.225 21.695 93.325 21.700 ;
        RECT 120.205 21.695 121.305 21.700 ;
        RECT 61.925 21.445 64.030 21.695 ;
        RECT 88.920 21.445 91.025 21.695 ;
        RECT 92.215 21.445 94.320 21.695 ;
        RECT 119.210 21.445 121.315 21.695 ;
        RECT 61.935 21.440 63.035 21.445 ;
        RECT 89.915 21.440 91.015 21.445 ;
        RECT 92.225 21.440 93.325 21.445 ;
        RECT 120.205 21.440 121.305 21.445 ;
        RECT 121.760 21.050 126.505 22.155 ;
        RECT 60.390 20.660 126.505 21.050 ;
        RECT 60.390 19.560 61.285 20.660 ;
        RECT 61.935 20.215 63.035 20.220 ;
        RECT 89.915 20.215 91.015 20.220 ;
        RECT 92.225 20.215 93.325 20.220 ;
        RECT 120.205 20.215 121.305 20.220 ;
        RECT 61.925 19.965 64.030 20.215 ;
        RECT 88.920 19.965 91.025 20.215 ;
        RECT 92.215 19.965 94.320 20.215 ;
        RECT 119.210 19.965 121.315 20.215 ;
        RECT 61.935 19.960 63.035 19.965 ;
        RECT 89.915 19.960 91.015 19.965 ;
        RECT 92.225 19.960 93.325 19.965 ;
        RECT 120.205 19.960 121.305 19.965 ;
        RECT 121.760 19.560 126.505 20.660 ;
        RECT 60.390 19.170 126.505 19.560 ;
        RECT 60.390 18.110 61.285 19.170 ;
        RECT 61.935 18.735 63.035 18.740 ;
        RECT 89.920 18.735 91.020 18.740 ;
        RECT 92.225 18.735 93.325 18.740 ;
        RECT 120.205 18.735 121.305 18.740 ;
        RECT 61.925 18.485 64.030 18.735 ;
        RECT 88.920 18.485 91.025 18.735 ;
        RECT 92.215 18.485 94.320 18.735 ;
        RECT 119.210 18.485 121.315 18.735 ;
        RECT 61.935 18.480 63.035 18.485 ;
        RECT 89.920 18.480 91.020 18.485 ;
        RECT 92.225 18.480 93.325 18.485 ;
        RECT 120.205 18.480 121.305 18.485 ;
        RECT 121.760 18.110 126.505 19.170 ;
        RECT 60.390 17.720 126.505 18.110 ;
        RECT 126.940 18.030 127.190 19.075 ;
        RECT 60.390 16.640 61.285 17.720 ;
        RECT 61.935 17.255 63.035 17.260 ;
        RECT 89.915 17.255 91.015 17.260 ;
        RECT 92.225 17.255 93.325 17.260 ;
        RECT 120.205 17.255 121.305 17.260 ;
        RECT 61.925 17.005 64.030 17.255 ;
        RECT 88.920 17.005 91.025 17.255 ;
        RECT 92.215 17.005 94.320 17.255 ;
        RECT 119.210 17.005 121.315 17.255 ;
        RECT 61.935 17.000 63.035 17.005 ;
        RECT 89.915 17.000 91.015 17.005 ;
        RECT 92.225 17.000 93.325 17.005 ;
        RECT 120.205 17.000 121.305 17.005 ;
        RECT 121.760 16.640 126.505 17.720 ;
        RECT 126.885 17.030 127.245 18.030 ;
        RECT 126.940 16.970 127.190 17.030 ;
        RECT 60.340 16.490 126.535 16.640 ;
        RECT 127.690 16.490 128.040 41.495 ;
        RECT 128.420 41.010 128.670 41.070 ;
        RECT 128.365 40.010 128.725 41.010 ;
        RECT 128.420 38.965 128.670 40.010 ;
        RECT 128.420 18.030 128.670 19.075 ;
        RECT 128.365 17.030 128.725 18.030 ;
        RECT 128.420 16.970 128.670 17.030 ;
        RECT 129.100 16.490 129.450 41.495 ;
        RECT 129.900 41.010 130.150 41.070 ;
        RECT 129.845 40.010 130.205 41.010 ;
        RECT 129.900 38.965 130.150 40.010 ;
        RECT 129.900 18.030 130.150 19.075 ;
        RECT 129.845 17.030 130.205 18.030 ;
        RECT 129.900 16.970 130.150 17.030 ;
        RECT 130.590 16.490 130.940 41.495 ;
        RECT 131.380 41.010 131.630 41.070 ;
        RECT 131.325 40.010 131.685 41.010 ;
        RECT 131.380 38.965 131.630 40.010 ;
        RECT 131.380 18.030 131.630 19.075 ;
        RECT 131.325 17.030 131.685 18.030 ;
        RECT 131.380 16.970 131.630 17.030 ;
        RECT 132.085 16.490 132.435 41.495 ;
        RECT 132.860 41.010 133.110 41.070 ;
        RECT 132.805 40.010 133.165 41.010 ;
        RECT 132.860 38.965 133.110 40.010 ;
        RECT 133.620 27.055 134.480 41.495 ;
        RECT 137.560 28.680 137.880 28.740 ;
        RECT 137.540 28.335 137.900 28.680 ;
        RECT 137.560 28.275 137.880 28.335 ;
        RECT 133.620 26.395 136.850 27.055 ;
        RECT 132.860 18.030 133.110 19.075 ;
        RECT 132.805 17.030 133.165 18.030 ;
        RECT 132.860 16.970 133.110 17.030 ;
        RECT 133.620 16.490 134.795 26.395 ;
        RECT 135.295 26.005 135.545 26.065 ;
        RECT 135.240 25.005 135.600 26.005 ;
        RECT 135.295 23.960 135.545 25.005 ;
        RECT 135.295 18.025 135.545 19.070 ;
        RECT 135.240 17.025 135.600 18.025 ;
        RECT 135.295 16.965 135.545 17.025 ;
        RECT 136.060 16.555 136.770 26.395 ;
        RECT 135.900 16.490 136.790 16.555 ;
        RECT 60.340 15.635 136.790 16.490 ;
        RECT 137.550 16.170 138.020 16.230 ;
        RECT 137.530 15.720 138.040 16.170 ;
        RECT 137.550 15.660 138.020 15.720 ;
        RECT 125.670 15.585 136.790 15.635 ;
        RECT 135.900 15.555 136.790 15.585 ;
      LAYER met2 ;
        RECT 60.960 58.465 120.110 58.585 ;
        RECT 60.960 57.705 122.995 58.465 ;
        RECT 60.960 53.305 61.580 57.705 ;
        RECT 62.170 56.275 62.430 57.705 ;
        RECT 65.360 56.275 65.620 57.705 ;
        RECT 69.845 56.275 70.105 57.705 ;
        RECT 73.040 56.275 73.300 57.705 ;
        RECT 76.235 56.275 76.495 57.705 ;
        RECT 79.430 56.275 79.690 57.705 ;
        RECT 82.625 56.275 82.885 57.705 ;
        RECT 85.820 56.275 86.080 57.705 ;
        RECT 89.015 56.275 89.275 57.705 ;
        RECT 92.210 56.275 92.470 57.705 ;
        RECT 95.405 56.275 95.665 57.705 ;
        RECT 98.600 56.275 98.860 57.705 ;
        RECT 101.795 56.275 102.055 57.705 ;
        RECT 104.990 56.270 105.250 57.705 ;
        RECT 106.895 56.270 107.155 57.705 ;
        RECT 110.090 56.270 110.350 57.705 ;
        RECT 113.285 56.270 113.545 57.705 ;
        RECT 116.480 56.270 116.740 57.705 ;
        RECT 118.505 57.395 122.995 57.705 ;
        RECT 118.505 57.365 120.110 57.395 ;
        RECT 62.525 54.285 62.925 54.645 ;
        RECT 53.450 52.070 60.145 52.095 ;
        RECT 53.430 51.810 60.145 52.070 ;
        RECT 62.525 51.810 62.815 54.285 ;
        RECT 53.430 51.510 62.815 51.810 ;
        RECT 53.430 51.220 60.145 51.510 ;
        RECT 53.450 51.195 60.145 51.220 ;
        RECT 45.580 47.655 59.710 47.660 ;
        RECT 45.580 47.650 60.915 47.655 ;
        RECT 45.580 44.565 61.260 47.650 ;
        RECT 62.525 46.755 62.815 51.510 ;
        RECT 63.460 52.150 63.720 55.295 ;
        RECT 65.715 54.285 66.115 54.645 ;
        RECT 63.460 51.750 63.755 52.150 ;
        RECT 62.525 46.395 62.925 46.755 ;
        RECT 62.170 44.565 62.430 45.810 ;
        RECT 63.460 45.790 63.720 51.750 ;
        RECT 65.715 48.760 66.005 54.285 ;
        RECT 66.650 50.465 66.910 55.295 ;
        RECT 68.555 54.795 75.205 55.295 ;
        RECT 78.140 54.795 84.790 55.295 ;
        RECT 87.725 54.795 94.375 55.295 ;
        RECT 97.310 55.290 103.715 55.295 ;
        RECT 97.310 54.795 103.960 55.290 ;
        RECT 68.555 51.305 68.815 54.795 ;
        RECT 69.350 54.280 69.750 54.640 ;
        RECT 72.545 54.285 72.945 54.645 ;
        RECT 75.740 54.285 76.140 54.645 ;
        RECT 68.540 50.885 68.860 51.305 ;
        RECT 66.650 50.065 66.950 50.465 ;
        RECT 65.715 48.360 66.015 48.760 ;
        RECT 65.715 46.770 66.005 48.360 ;
        RECT 65.715 46.410 66.115 46.770 ;
        RECT 65.360 44.565 65.620 45.825 ;
        RECT 66.650 45.805 66.910 50.065 ;
        RECT 68.555 45.805 68.815 50.885 ;
        RECT 69.460 46.770 69.750 54.280 ;
        RECT 72.655 46.770 72.945 54.285 ;
        RECT 75.850 53.955 76.140 54.285 ;
        RECT 75.780 53.300 76.265 53.955 ;
        RECT 75.850 46.770 76.140 53.300 ;
        RECT 78.140 49.625 78.400 54.795 ;
        RECT 78.935 54.285 79.335 54.645 ;
        RECT 82.130 54.285 82.530 54.645 ;
        RECT 85.325 54.285 85.725 54.645 ;
        RECT 78.105 49.190 78.440 49.625 ;
        RECT 69.350 46.410 69.750 46.770 ;
        RECT 72.545 46.410 72.945 46.770 ;
        RECT 75.740 46.410 76.140 46.770 ;
        RECT 78.140 45.805 78.400 49.190 ;
        RECT 79.045 46.770 79.335 54.285 ;
        RECT 82.240 46.770 82.530 54.285 ;
        RECT 85.435 54.005 85.725 54.285 ;
        RECT 85.370 53.350 85.855 54.005 ;
        RECT 85.435 46.770 85.725 53.350 ;
        RECT 78.935 46.410 79.335 46.770 ;
        RECT 82.130 46.410 82.530 46.770 ;
        RECT 85.325 46.410 85.725 46.770 ;
        RECT 87.725 52.245 87.985 54.795 ;
        RECT 88.520 54.285 88.920 54.645 ;
        RECT 91.715 54.285 92.115 54.645 ;
        RECT 94.910 54.285 95.310 54.645 ;
        RECT 87.725 51.845 88.025 52.245 ;
        RECT 87.725 45.805 87.985 51.845 ;
        RECT 88.630 46.770 88.920 54.285 ;
        RECT 91.825 46.770 92.115 54.285 ;
        RECT 95.020 53.970 95.310 54.285 ;
        RECT 94.905 53.315 95.390 53.970 ;
        RECT 95.020 46.770 95.310 53.315 ;
        RECT 88.520 46.410 88.920 46.770 ;
        RECT 91.715 46.410 92.115 46.770 ;
        RECT 94.910 46.410 95.310 46.770 ;
        RECT 97.310 50.455 97.570 54.795 ;
        RECT 103.700 54.790 103.960 54.795 ;
        RECT 101.410 54.645 101.700 54.655 ;
        RECT 98.105 54.285 98.505 54.645 ;
        RECT 101.300 54.285 101.700 54.645 ;
        RECT 104.605 54.640 104.895 54.650 ;
        RECT 97.310 50.005 97.660 50.455 ;
        RECT 97.310 45.805 97.570 50.005 ;
        RECT 98.215 46.770 98.505 54.285 ;
        RECT 101.410 46.770 101.700 54.285 ;
        RECT 104.495 54.280 104.895 54.640 ;
        RECT 104.605 53.990 104.895 54.280 ;
        RECT 107.250 54.640 107.540 54.730 ;
        RECT 107.250 54.280 107.650 54.640 ;
        RECT 104.530 53.335 105.015 53.990 ;
        RECT 104.605 46.770 104.895 53.335 ;
        RECT 107.250 51.310 107.540 54.280 ;
        RECT 107.235 50.875 107.555 51.310 ;
        RECT 98.105 46.410 98.505 46.770 ;
        RECT 101.300 46.410 101.700 46.770 ;
        RECT 104.495 46.410 104.895 46.770 ;
        RECT 107.250 46.770 107.540 50.875 ;
        RECT 108.185 48.250 108.445 55.290 ;
        RECT 110.445 54.640 110.735 54.770 ;
        RECT 110.445 54.280 110.845 54.640 ;
        RECT 110.445 49.630 110.735 54.280 ;
        RECT 111.380 49.640 111.640 55.290 ;
        RECT 113.640 54.640 113.930 54.755 ;
        RECT 113.640 54.280 114.040 54.640 ;
        RECT 113.640 52.270 113.930 54.280 ;
        RECT 113.640 51.820 113.950 52.270 ;
        RECT 110.415 49.180 110.825 49.630 ;
        RECT 111.380 49.190 111.730 49.640 ;
        RECT 108.185 47.850 108.485 48.250 ;
        RECT 107.250 46.410 107.650 46.770 ;
        RECT 67.140 44.565 68.000 44.590 ;
        RECT 45.580 44.375 68.000 44.565 ;
        RECT 106.895 44.520 107.155 45.825 ;
        RECT 108.185 45.805 108.445 47.850 ;
        RECT 110.445 46.770 110.735 49.180 ;
        RECT 110.445 46.410 110.845 46.770 ;
        RECT 110.090 44.520 110.350 45.825 ;
        RECT 111.380 45.805 111.640 49.190 ;
        RECT 113.640 46.770 113.930 51.820 ;
        RECT 114.575 51.705 114.835 55.290 ;
        RECT 116.835 54.640 117.125 54.775 ;
        RECT 116.835 54.280 117.235 54.640 ;
        RECT 114.575 51.205 114.975 51.705 ;
        RECT 113.640 46.410 114.040 46.770 ;
        RECT 113.285 44.520 113.545 45.825 ;
        RECT 114.575 45.805 114.835 51.205 ;
        RECT 116.835 50.480 117.125 54.280 ;
        RECT 117.770 52.740 118.030 55.290 ;
        RECT 118.505 53.360 119.125 57.365 ;
        RECT 117.770 52.290 129.915 52.740 ;
        RECT 116.835 49.980 117.170 50.480 ;
        RECT 116.835 46.770 117.125 49.980 ;
        RECT 116.835 46.410 117.235 46.770 ;
        RECT 116.480 44.520 116.740 45.825 ;
        RECT 117.770 45.805 118.030 52.290 ;
        RECT 120.030 46.770 120.330 48.275 ;
        RECT 123.225 46.770 123.525 49.665 ;
        RECT 126.420 46.770 126.720 51.730 ;
        RECT 129.615 46.770 129.915 52.290 ;
        RECT 120.030 46.410 120.430 46.770 ;
        RECT 123.225 46.410 123.625 46.770 ;
        RECT 126.420 46.410 126.820 46.770 ;
        RECT 129.615 46.410 130.015 46.770 ;
        RECT 126.065 44.545 126.325 45.925 ;
        RECT 125.380 44.520 126.890 44.545 ;
        RECT 106.400 44.475 119.200 44.520 ;
        RECT 45.580 44.370 59.710 44.375 ;
        RECT 60.420 43.605 68.000 44.375 ;
        RECT 60.420 43.270 61.260 43.605 ;
        RECT 67.140 42.685 68.000 43.605 ;
        RECT 69.845 43.325 72.010 43.825 ;
        RECT 73.040 43.325 75.205 43.825 ;
        RECT 76.235 42.685 76.495 43.825 ;
        RECT 79.430 43.325 81.595 43.825 ;
        RECT 82.625 43.325 84.790 43.825 ;
        RECT 85.820 42.685 86.080 43.825 ;
        RECT 89.015 43.325 91.180 43.825 ;
        RECT 92.210 43.325 94.375 43.825 ;
        RECT 95.405 43.395 95.665 43.825 ;
        RECT 95.405 43.325 95.670 43.395 ;
        RECT 98.600 43.325 100.765 43.825 ;
        RECT 101.795 43.325 103.960 43.825 ;
        RECT 95.410 42.685 95.670 43.325 ;
        RECT 104.990 42.685 105.250 43.825 ;
        RECT 105.750 43.465 119.200 44.475 ;
        RECT 105.750 42.685 106.815 43.465 ;
        RECT 67.140 41.630 106.815 42.685 ;
        RECT 67.140 41.610 106.145 41.630 ;
        RECT 56.990 19.350 57.890 39.135 ;
        RECT 118.455 35.645 119.200 43.465 ;
        RECT 124.915 43.840 126.890 44.520 ;
        RECT 124.915 42.005 125.470 43.840 ;
        RECT 127.355 42.665 127.615 45.925 ;
        RECT 129.260 44.565 129.520 45.925 ;
        RECT 128.050 43.860 129.860 44.565 ;
        RECT 130.550 43.505 130.810 45.925 ;
        RECT 130.550 43.245 137.850 43.505 ;
        RECT 127.355 42.405 135.550 42.665 ;
        RECT 119.675 35.645 119.935 41.425 ;
        RECT 118.455 34.895 120.265 35.645 ;
        RECT 120.965 30.630 121.255 41.425 ;
        RECT 122.870 35.620 123.130 41.425 ;
        RECT 124.160 41.060 127.195 41.425 ;
        RECT 124.160 36.325 124.420 41.060 ;
        RECT 124.935 35.620 125.495 40.755 ;
        RECT 126.935 39.960 127.195 41.060 ;
        RECT 128.415 40.700 130.155 41.060 ;
        RECT 128.415 39.960 128.675 40.700 ;
        RECT 129.895 39.960 130.155 40.700 ;
        RECT 131.375 40.700 133.115 41.060 ;
        RECT 131.375 39.960 131.635 40.700 ;
        RECT 132.855 39.960 133.115 40.700 ;
        RECT 121.800 34.850 125.495 35.620 ;
        RECT 61.985 30.270 62.985 30.630 ;
        RECT 89.965 30.270 93.275 30.630 ;
        RECT 120.255 30.270 121.255 30.630 ;
        RECT 61.985 29.150 62.345 30.270 ;
        RECT 61.985 28.790 62.985 29.150 ;
        RECT 89.965 28.790 93.275 29.150 ;
        RECT 120.255 28.790 121.255 29.150 ;
        RECT 120.895 27.670 121.255 28.790 ;
        RECT 61.985 27.310 62.985 27.670 ;
        RECT 89.965 27.310 93.275 27.670 ;
        RECT 120.255 27.310 121.255 27.670 ;
        RECT 61.985 26.190 62.345 27.310 ;
        RECT 61.985 25.830 62.985 26.190 ;
        RECT 89.965 25.830 93.275 26.190 ;
        RECT 120.255 25.830 121.255 26.190 ;
        RECT 120.895 24.710 121.255 25.830 ;
        RECT 135.290 24.955 135.550 42.405 ;
        RECT 137.590 28.285 137.850 43.245 ;
        RECT 61.985 24.350 62.985 24.710 ;
        RECT 89.965 24.350 93.275 24.710 ;
        RECT 120.255 24.350 121.255 24.710 ;
        RECT 61.985 23.230 62.345 24.350 ;
        RECT 61.985 22.870 62.985 23.230 ;
        RECT 89.965 22.870 93.275 23.230 ;
        RECT 120.255 22.870 121.255 23.230 ;
        RECT 120.895 21.750 121.255 22.870 ;
        RECT 61.985 21.390 62.985 21.750 ;
        RECT 89.965 21.390 93.275 21.750 ;
        RECT 120.255 21.390 121.255 21.750 ;
        RECT 61.985 20.270 62.345 21.390 ;
        RECT 61.985 19.910 62.985 20.270 ;
        RECT 89.965 19.910 93.275 20.270 ;
        RECT 120.255 19.910 121.255 20.270 ;
        RECT 56.970 18.500 57.910 19.350 ;
        RECT 120.895 18.790 121.255 19.910 ;
        RECT 56.990 18.475 57.890 18.500 ;
        RECT 61.985 18.430 62.985 18.790 ;
        RECT 89.970 18.430 93.275 18.790 ;
        RECT 120.255 18.430 121.255 18.790 ;
        RECT 61.985 17.310 62.345 18.430 ;
        RECT 126.935 17.340 127.195 18.080 ;
        RECT 128.415 17.340 128.675 18.080 ;
        RECT 61.985 16.950 62.985 17.310 ;
        RECT 89.965 16.950 93.275 17.310 ;
        RECT 120.255 16.950 124.030 17.310 ;
        RECT 126.935 16.980 128.675 17.340 ;
        RECT 129.895 17.340 130.155 18.080 ;
        RECT 131.375 17.340 131.635 18.080 ;
        RECT 129.895 16.980 131.635 17.340 ;
        RECT 123.670 15.395 124.030 16.950 ;
        RECT 132.855 15.395 133.115 18.080 ;
        RECT 135.290 15.395 135.550 18.075 ;
        RECT 137.580 15.395 137.990 16.220 ;
        RECT 123.670 15.035 137.990 15.395 ;
        RECT 136.170 9.310 137.070 15.035 ;
        RECT 136.150 8.460 137.090 9.310 ;
        RECT 136.170 8.435 137.070 8.460 ;
      LAYER met3 ;
        RECT 121.905 58.465 122.975 58.490 ;
        RECT 121.905 57.395 129.715 58.465 ;
        RECT 121.905 57.370 122.975 57.395 ;
        RECT 62.475 53.165 62.865 53.190 ;
        RECT 91.775 53.165 92.165 53.190 ;
        RECT 101.360 53.165 101.750 53.190 ;
        RECT 62.475 52.865 101.895 53.165 ;
        RECT 62.475 52.840 62.865 52.865 ;
        RECT 91.775 52.840 92.165 52.865 ;
        RECT 101.360 52.840 101.750 52.865 ;
        RECT 113.590 52.220 114.000 52.245 ;
        RECT 63.410 52.100 63.805 52.125 ;
        RECT 72.605 52.100 72.995 52.125 ;
        RECT 82.190 52.100 82.580 52.125 ;
        RECT 53.450 48.470 54.350 52.095 ;
        RECT 63.410 51.800 82.760 52.100 ;
        RECT 87.675 51.870 114.000 52.220 ;
        RECT 113.590 51.845 114.000 51.870 ;
        RECT 63.410 51.775 63.805 51.800 ;
        RECT 72.605 51.775 72.995 51.800 ;
        RECT 82.190 51.775 82.580 51.800 ;
        RECT 126.370 51.680 126.770 51.705 ;
        RECT 68.490 50.910 69.315 51.280 ;
        RECT 106.925 50.900 107.605 51.285 ;
        RECT 114.525 51.230 126.770 51.680 ;
        RECT 126.370 51.205 126.770 51.230 ;
        RECT 66.600 50.415 67.000 50.440 ;
        RECT 69.410 50.415 69.800 50.440 ;
        RECT 88.580 50.415 88.970 50.440 ;
        RECT 116.785 50.430 117.220 50.455 ;
        RECT 66.600 50.115 89.025 50.415 ;
        RECT 66.600 50.090 67.000 50.115 ;
        RECT 69.410 50.090 69.800 50.115 ;
        RECT 88.580 50.090 88.970 50.115 ;
        RECT 97.260 50.030 117.220 50.430 ;
        RECT 116.785 50.005 117.220 50.030 ;
        RECT 123.175 49.615 123.575 49.640 ;
        RECT 78.055 49.215 78.990 49.600 ;
        RECT 109.950 49.205 110.875 49.605 ;
        RECT 111.330 49.215 123.575 49.615 ;
        RECT 123.175 49.190 123.575 49.215 ;
        RECT 65.665 48.710 66.065 48.735 ;
        RECT 78.995 48.710 79.385 48.735 ;
        RECT 98.165 48.710 98.555 48.735 ;
        RECT 53.455 48.445 54.345 48.470 ;
        RECT 65.665 48.410 101.895 48.710 ;
        RECT 65.665 48.385 66.065 48.410 ;
        RECT 78.995 48.385 79.385 48.410 ;
        RECT 98.165 48.385 98.555 48.410 ;
        RECT 119.980 48.225 120.380 48.250 ;
        RECT 108.135 47.875 120.380 48.225 ;
        RECT 119.980 47.850 120.380 47.875 ;
        RECT 45.600 47.660 48.890 47.685 ;
        RECT 35.590 44.370 48.890 47.660 ;
        RECT 45.600 44.345 48.890 44.370 ;
        RECT 56.990 12.365 57.890 19.375 ;
        RECT 56.965 11.475 57.915 12.365 ;
        RECT 56.990 11.470 57.890 11.475 ;
        RECT 136.170 6.195 137.070 9.335 ;
        RECT 136.145 5.305 137.095 6.195 ;
        RECT 136.170 5.300 137.070 5.305 ;
      LAYER met4 ;
        RECT 15.025 224.760 15.030 224.935 ;
        RECT 17.785 224.760 17.790 224.870 ;
        RECT 20.850 224.760 20.855 224.905 ;
        RECT 15.025 220.545 15.330 224.760 ;
        RECT 17.785 220.545 18.090 224.760 ;
        RECT 20.550 220.545 20.855 224.760 ;
        RECT 23.305 224.760 23.310 224.895 ;
        RECT 26.370 224.760 26.375 224.945 ;
        RECT 29.130 224.760 29.135 224.895 ;
        RECT 23.305 220.545 23.610 224.760 ;
        RECT 26.070 220.545 26.375 224.760 ;
        RECT 28.830 220.545 29.135 224.760 ;
        RECT 31.585 224.760 31.590 224.935 ;
        RECT 34.650 224.760 34.655 224.850 ;
        RECT 37.410 224.760 37.415 224.835 ;
        RECT 40.170 224.760 40.175 224.915 ;
        RECT 42.930 224.760 42.935 224.905 ;
        RECT 31.585 220.545 31.890 224.760 ;
        RECT 34.350 220.545 34.655 224.760 ;
        RECT 37.110 220.545 37.415 224.760 ;
        RECT 39.870 220.545 40.175 224.760 ;
        RECT 42.630 220.545 42.935 224.760 ;
        RECT 45.385 224.760 45.390 224.915 ;
        RECT 48.145 224.760 48.150 224.795 ;
        RECT 51.210 224.760 51.215 224.850 ;
        RECT 53.970 224.760 53.975 224.960 ;
        RECT 56.730 224.760 56.735 224.960 ;
        RECT 59.490 224.760 59.495 224.885 ;
        RECT 45.385 220.545 45.690 224.760 ;
        RECT 48.145 220.545 48.450 224.760 ;
        RECT 50.910 220.545 51.215 224.760 ;
        RECT 53.670 220.545 53.975 224.760 ;
        RECT 56.430 220.545 56.735 224.760 ;
        RECT 59.190 220.545 59.495 224.760 ;
        RECT 61.945 224.760 61.950 224.840 ;
        RECT 64.705 224.760 64.710 224.975 ;
        RECT 67.770 224.760 67.775 224.915 ;
        RECT 61.945 220.545 62.250 224.760 ;
        RECT 64.705 220.545 65.010 224.760 ;
        RECT 67.470 220.545 67.775 224.760 ;
        RECT 70.225 224.760 70.230 224.945 ;
        RECT 76.050 224.760 76.060 224.980 ;
        RECT 70.225 220.545 70.530 224.760 ;
        RECT 72.990 220.545 73.290 224.760 ;
        RECT 75.750 220.545 76.060 224.760 ;
        RECT 78.500 224.760 78.510 224.840 ;
        RECT 78.500 220.545 78.810 224.760 ;
        RECT 6.000 218.775 79.195 220.545 ;
        RECT 128.620 58.465 129.690 58.470 ;
        RECT 128.620 57.395 142.000 58.465 ;
        RECT 128.620 57.390 129.690 57.395 ;
        RECT 107.230 51.260 107.560 51.265 ;
        RECT 68.535 50.925 107.560 51.260 ;
        RECT 107.230 50.920 107.560 50.925 ;
        RECT 110.410 49.580 110.830 49.585 ;
        RECT 35.615 47.660 38.905 47.665 ;
        RECT 6.000 44.370 38.905 47.660 ;
        RECT 35.615 44.365 38.905 44.370 ;
        RECT 53.450 8.230 54.350 49.370 ;
        RECT 78.100 49.230 110.830 49.580 ;
        RECT 110.410 49.225 110.830 49.230 ;
        RECT 56.990 11.470 117.750 12.370 ;
        RECT 53.450 7.330 98.430 8.230 ;
        RECT 97.530 1.000 98.430 7.330 ;
        RECT 116.850 1.000 117.750 11.470 ;
        RECT 136.170 1.000 137.070 6.200 ;
  END
END tt_um_DalinEM_G_Control
END LIBRARY

